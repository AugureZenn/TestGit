test de fichier 
xcvcvxvxv